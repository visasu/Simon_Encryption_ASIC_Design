//NumStages defines the number of pipeline stages in Your design. Minimum Numstags = 1 is for non-pipelined design 
//i.e. no intermediate flip-flops between I/O flipflops.
localparam NumStages = 32;
// clock period in ns (nano second)
localparam ClkPeriod = 0.442;
